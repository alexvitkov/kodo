fn foo(x: i32) {};
fn foo(x: i16) {};
fn foo(x: u8) {};
fn foo(x: u16) {};
