fn foo() {};
fn foo(x: i32) {};
fn foo(x: i32, y: i32) {};
