fn foo(x: u32, y: u32) { };

a: u32;
b: u32;

foo(a, b); // this must find the global variables
