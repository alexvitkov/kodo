fn foo(x: i32) { };

x; // this must fail to resolve
