// functions cannot be overloaded by return type alone
fn foo(x: i32): i32 { };
fn foo(x: i32): u32 { };
