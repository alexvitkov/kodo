if (foo) { };

if (foo) { } else { };
