fn foo(x: i64) { };

x := 12345; // number_literal gets casted to i64 by default

foo(x);
