
fn foo[X] (x: X) {};
fn foo[X, Y] () {};
fn foo[X, Y, Z] () {};
