fn foo(x: i32, y: i32): u32 {};
fn foo(x: i32, y: i32): u32 {};
