x: i32;
y: u8;

fn foo[T1, T2](a: T1, b: T2) { };

foo(x, y);
