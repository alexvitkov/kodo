// make sure the := syntax works with a space in the middle
{ foo : = bar; };
{ foo := bar; };
