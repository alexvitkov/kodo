foo: i32;
foo: u16;
