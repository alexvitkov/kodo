fn foo(x) { }
