foo: i32;
foo: i32;
