// variables can be declared in the condition
// they must be available in then/else blocks
 
if (x: i32) {
    x;
} else {
    x;
};
