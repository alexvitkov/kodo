100;
0;
1000000000000000000000000000000000;
