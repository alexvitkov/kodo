foo();

foo(x, y, z);

foo(bar(), x, y, z);
