x: i32;
y := x; // y: i32

fn foo(x: i32, y: i32) { };

foo(x, y);
