// trailing comma is not allowed
fn foo(x: i32, ) { };
