{ a + (b * c); };
{ a + (b * c); };
