foo1: i8  = 100;
foo2: i32 = 100;
foo3: i64 = 100;
foo4: i64 = 100;
foo5: u8  = 100;
foo6: u32 = 100;
foo7: u64 = 100;
foo8: u64 = 100;
