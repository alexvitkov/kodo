x: i32;
y: i32;

fn foo[T](a: T, b: T) {};

foo(x, y);
