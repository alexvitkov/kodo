foo1: i8  = bar1: i8;
foo2: i16 = bar2: i16;
foo3: i32 = bar3: i32;
foo4: i64 = bar4: i64;
foo5: u8  = bar5: u8;
foo6: u16 = bar6: u16;
foo7: u32 = bar7: u32;
foo8: u64 = bar8: u64;
