fn foo(x: i32, y: i32) {
    foo(x, y); // this must find the arguments
};
