{
};

{
    ;
    ;
    ;
}

{
    foo();
    bar();
    baz();
};
