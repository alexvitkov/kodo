// empty block
{
};

// make sure empty expressions are allowed
{
    ;
    ;
    ;
}

// block with some elements
{
    foo();
    bar();
    baz();
};
