fn foo() {};
fn foo() {};
