fn () { };
fn foo() { };

fn (): i32 { };
fn bar(): i32 { };

fn (x: i32): i32 { };
fn baz(x: i32): i32 { };

fn (x: i32, y: i32): i32 { };
fn baz(x: i32, y: i32): i32 { };
